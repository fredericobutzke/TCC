
module inv ( A, Z )

(* integer foreign      = "SystemC";
*);
  input A;
  output Z;
endmodule
