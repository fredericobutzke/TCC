
module nand2 ( A, B, Z )

(* integer foreign      = "SystemC";
*);
  input A, B;
  output Z;
endmodule
